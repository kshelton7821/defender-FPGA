library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package data_etc is
	type game_entity is
	record
		entity_type : STD_LOGIC_VECTOR(2 downto 0);
		posx		: integer;
		posy		: integer;
		len			: integer;
		height		: integer;
		imageID 	: integer;
		enable 	: STD_LOGIC;
		toDelete : std_logic;
		expCount : integer range 0 to 500;
	end record;
	type entities is array (20 downto 0) of game_entity;
	constant playerPixels : STD_LOGIC_VECTOR(2499 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000001111111111111100000000000000000000000000000000111111111111111110000000000000000000000000000000001111111111111111100000000000000000000000000000011111111111111111000000000000000000000000000000000111111111111111110000000000000000000000000000000011111111111111111100000000000000000000000000000001111111111111111110000000000000000000000000000000011111111011111111000000000000000000000000000000001111111111111111110000000000000000000000000000011111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000011111111111111111110000000000000000000000001110111111111111111111111100000000000000000000000011101111111111101111111111000000000000000000000000011111111111111111111111110000000000000000111111111111111111111111111111111000000000000000001111111111111111111110000000000000000000000000000111111111111111111111111111111111100000000000000111111111111111110111111111111111111001111000000001111111111111111101111111111111111110011111100000110000111111000000111111110000000000000111111000011111111111111111111111111111111111111001111111000111111110111111111111111111111111111110011111110001111111101111111111111111111111111111100111111100011111111111111111111111111111111111111001111111000011000011111100000011111111000000000000011111100000011111111111111111011111111111111111100111111000000111111111111111110111111111111111111001111000000000011111111111111111111111111111111110000000000000000011111111111111111111100000000000000000000000000000111111111111111111111111111111111000000000000000000000000001111111111111111111111111000000000000000000000000111011111111111011111111110000000000000000000000001110111111111111111111111100000000000000000000000000000001111111111111111111000000000000000000000000000000001111111111000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000111111111111111111000000000000000000000000000000000111111110111111110000000000000000000000000000000001111111111111111110000000000000000000000000000000001111111111111111110000000000000000000000000000000001111111111111111100000000000000000000000000000000011111111111111111000000000000000000000000000000000000111111111111111110000000000000000000000000000000001111111111111111100000000000000000000000000000000000001111111111111100000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000";
	constant alien1Pixels : STD_LOGIC_VECTOR(2499 downto 0) := "0000000000000111111111111100000000001111111111111100000000000001111111111111000000000011111111111111000000000000011111111111110000000000111111111111100000000000000111111111111100000000001111111111111000000000000001111111111111000011111111111111111110000000000000011111111111110000111111111111111111100000000000000111111011111100001111111111111111111000000000000011111110111111000011111111111111111110000000000001111111101111110000111111111111111111110000000000011111111011111100001111111111111111111100000000000111111110111111000011111111111111111110000000000001111111101111110000111111111111100000000000000000001111111011111100001111111111111000000000000000000000011110111111000011111111111110000000000000000000011111111111111111111111111111100000000000000000000111111111111111111111111100000000000000000000000001111111111111111111111111100000000000000000000000011111111111111111111111110000000000000111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111100000000000000111111111111111111111111111111111111000000000000001111111111111111111111111111111111110000000000000111111111111111111111111111111111111100111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111110000000000000000001011111111111111111111111110000000000000000000000000111111111111111111111111100000000000000000000000001111111111111111111111111010000000000000000000000011111111111111111111111111111100000000000000000000111111011111111111111111111111000000000000000000011111110111111000011111111111110000000000000000001111111101111110000111111111111100000000000000000011111111011111100001111111111111111111000000000000111111110111111000011111111111111111110000000000001111111101111110000111111111111111111110000000000001111111011111100001111111111111111111000000000000000011110111111000011111111111111111110000000000000011111111111110000111111111111111111100000000000000111111111111100001111111111111111111000000000000001111111111111000000000011111111111110000000000000011111111111110000000000111111111111100000000000000111111111111100000000001111111111111000000000000001111111111111000000000011111111111101";
	constant alien2Pixels : STD_LOGIC_VECTOR(5999 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111101001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000111111011111111000000000000000000000000000000000001101111111111111111111111111111111111111111111111100000000000000000000000000000000000000000111101111111111111111101111100001111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000001111101111101111111111111111110111111111111111100000000000000000111111111111111111111111111111111111111111111111111111110110000000000000000000000000011111111000111111111111111111111100111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000001110011111111111111111111111111111111111111111111111111111000000000001100111111111111111111111111111111111111111111111111111111111110000000000000000011111111111011111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111011111111110000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111100111111111111111110000000011111011111111111111100001111111111111111111111111111110000111111111111111111111111000000000000000000000000000111110010010000000000001111111111111111111111001111111111111111111111111111111111111111111111111111111111111011100011111111110011100000000000000000000011100000011000000011111111111111111111111111000111111111111111111110111111111111111111111111111111111111111111111111111111111111111111000000000000000001000001100001111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000010111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000110111111111111111111111111111111111111111110000000000000000000011111111111111111111111111100110111100001111111111111111111111111100000000000000000001100011111111111111111111111111111111111111110000000000000000000000011111111111111111111111101111111100000000111111111111111111000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000011111111111111111111111101111111111111111110000000000000001110000000000000000001110000111111111111111111111111111111111111111000000000000000000000000011111111111111111111111101111111111111111111111111111000000111110000000000001111000011111111111111111111111111111111111111110000000000000000000000000000011111111111111111111000111111111111111111111111111111000011111111011111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111111111000000011111111111111111111111111111001111111010111101011111111111111111111111111111111111111111111000000000000000000000000000000000000001111111111110000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000111100000000000000000000001111111111111111111111111111111111111111110111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	constant alien3Pixels : STD_LOGIC_VECTOR(2799 downto 0) := "0000000111111111111111111111111110000000000000000000000001111111111111111111111111110000000000000000000000011111111111111111111111111110000000000000000000001111111111111111111111111111111100000000000000000011111111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000001111111111111111111111111111111110010000000000000011111111111111111111111111111111111100000000000000111111111111111111111111111111111111000000000000001111111111111111111111111111111111110000000000000001111111111111111111111111111111111100000000000000000000011111111111111111111111111110000000000000000000000111111111111111111111111111100000000000000000000011111111111111111111111111111110000000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111100000000000111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111100000000000001111111111111111111111111111111111110000000000000011111111111111111111111111111111110000000000000000001011111111111111111111111111111000000000000000000001011111111111111111111111111000000000000000000000011111111111111111111111111000000000000000000111111111111111111111111111111111110000000000000011111111111111111111111111111111111100000000000000111111111111111111111111111111111101000000000000011111111111111111111111111111111111110000000000000011111111111111111111111111111111111100000000000000111111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000000011111111111111111111111111111111000000000000000000011111111111111111111111111110000000000000000000000111111111111111111111111111000000000000000000000001111111111111111111111111100000000000000000";
	constant asteroidPixels : STD_LOGIC_VECTOR(3599 downto 0) := "000000000000000000000001110000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111000000000011111011111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111100000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000111100111111000000000000000000000000000000000000000000000000000000011000000000000000000000000000";
	constant explosionPixels : STD_LOGIC_VECTOR(2499 downto 0) := "0000000000000000000011000000110000000000000000000000000000000000000111111101111111100000000000000000000000000000000111111111111111111110000000000000000000000000000111111111111111111111111000000000000000000000000011111111111111111111111111000000000000000000000011111111111111111111111111111100000000000000000001111111111111111111111111111111100000000000000000111111111111111111111111111111111100000000000000011111111111111111111111111111111111100000000000001111111111111111111111111111111111111100000000000111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111110000001111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111000000000011111111111111111111111111111111111111110000000000011111111111111111111111111111111111111000000000000011111111111111111111111111111111111100000000000000011111111111111111111111111111111110000000000000000011111111111111111111111111111111000000000000000000011111111111111111111111111111100000000000000000000001111111111111111111111111100000000000000000000000001111111111111111111111110000000000000000000000000000111111111111111111110000000000000000000000000000000001111111111111100000000000000000000000000000000000000001111110000000000000000000000";
end package data_etc;